/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  ram_fball_down
(
		input [8:0] read_address,
		output logic [23:0] output_color
);

// mem has width of 3 bits and a total of 400 addresses
logic [3:0] mem [0:440];

logic [23:0] pal [3:0];
assign pal[0] = 24'h800080;
assign pal[1] = 24'hFFFFFF;
assign pal[2] = 24'hF83800;
assign pal[3] = 24'hFFA044;

assign output_color = pal[mem[read_address]];

initial
begin
	 $readmemh("C:/ece385/final_project/ECE385-HelperTools-master/PNG To Hex/On-Chip Memory/sprite_bytes/fball_down.txt", mem);
end

endmodule
