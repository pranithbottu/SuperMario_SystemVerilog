/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  ram_qblock_blink_2
(
		input [8:0] read_address,
		output logic [23:0] output_color
);

// mem has width of 4 bits and a total of 400 addresses
logic [3:0] mem [0:399];

logic [23:0] pal [4:0];
assign pal[0] = 24'h800080;
assign pal[1] = 24'h000000;
assign pal[2] = 24'hE75A10;
assign pal[3] = 24'hFFA542;
assign pal[4] = 24'h8C1000;

assign output_color = pal[mem[read_address]];

initial
begin
	 $readmemh("C:/ece385/final_project/ECE385-HelperTools-master/PNG To Hex/On-Chip Memory/sprite_bytes/qblock_blink_2.txt", mem);
end

endmodule
